----------------------------------------------------------------------------
-- Entity:        LightShowROM
-- Written By:    Robert Myers
-- Date Created:  11 Apr 22
-- Description:   VHDL model of a hex digit to 7-segment display ROM
--
-- Revision History (date, initials, description):
--
-- Dependencies:
--   (none)
----------------------------------------------------------------------------
library IEEE;
use     IEEE.STD_LOGIC_1164.ALL;
use     IEEE.NUMERIC_STD.ALL;

----------------------------------------------------------------------------
entity LightShowROM is
    port (
        A  : in  STD_LOGIC_VECTOR(7 downto 0);
        RD : out STD_LOGIC_VECTOR(31 downto 0)
    );
end entity;
----------------------------------------------------------------------------

architecture Behavioral of LightShowROM is

	type ROM_TYPE is ARRAY (0 to 255) of STD_LOGIC_VECTOR(31 downto 0);
	constant ROM : ROM_TYPE := (
	--  4-digit   LEDs                
		x"1000" & "1000000000000001", -- Address =   0
		x"0100" & "0100000000000010", -- Address =   1
		x"0010" & "0010000000000100", -- Address =   2
		x"0001" & "0001000000001000", -- Address =   3
		x"0002" & "0000100000010000", -- Address =   4
		x"0007" & "0000010000100000", -- Address =   5
		x"0070" & "0000001001000000", -- Address =   6
		x"0700" & "0000000110000000", -- Address =   7
		x"7000" & "0000000110000000", -- Address =   8
		x"5000" & "0000001001000000", -- Address =   9
		x"4000" & "0000010000100000", -- Address =  10
		x"0400" & "0000100000010000", -- Address =  11
		x"0040" & "0001000000001000", -- Address =  12
		x"0004" & "0010000000000100", -- Address =  13
		x"0003" & "0100000000000010", -- Address =  14
		x"0007" & "1000000000000001", -- Address =  15
		x"0070" & "1100000000000011", -- Address =  16
		x"0700" & "0110000000000110", -- Address =  17
		x"7000" & "0011000000001100", -- Address =  18
		x"0008" & "0001100000011000", -- Address =  19
		x"0089" & "0000110000110000", -- Address =  20
		x"089A" & "0000011001100000", -- Address =  21
		x"89AB" & "0000001111000000", -- Address =  22
		x"9ABC" & "0000000110000000", -- Address =  23
		x"ABC0" & "0000001111000000", -- Address =  24
		x"BC0D" & "0000011001100000", -- Address =  25
		x"C0DE" & "0000110000110000", -- Address =  26
		x"0DEF" & "0001100000011000", -- Address =  27
		x"DEF0" & "0011000000001100", -- Address =  28
		x"EF00" & "0110000000000110", -- Address =  29
		x"F000" & "1100000000000011", -- Address =  30
		x"0000" & "1110000000000111", -- Address =  31
		x"1100" & "0111000000001110", -- Address =  32
		x"0044" & "0011100000011100", -- Address =  33
		x"0011" & "0001110000111000", -- Address =  34
		x"4400" & "0000111001110000", -- Address =  35
		x"4141" & "0000011111100000", -- Address =  36
		x"1414" & "0000001111000000", -- Address =  37
		x"4141" & "0000001111000000", -- Address =  38
		x"1414" & "0000011111100000", -- Address =  39
		x"1000" & "0000111001110000", -- Address =  40
		x"0700" & "0001110000111000", -- Address =  41
		x"0040" & "0011100000011100", -- Address =  42
		x"0007" & "0111000000001110", -- Address =  43
		x"0010" & "1110000000000111", -- Address =  44
		x"0700" & "1111000000001111", -- Address =  45
		x"4000" & "0111100000011110", -- Address =  46
		x"0100" & "0011110000111100", -- Address =  47
		x"0010" & "0001111001111000", -- Address =  48
		x"0001" & "0000111111110000", -- Address =  49
		x"0002" & "0000011111100000", -- Address =  50
		x"0003" & "0000001111000000", -- Address =  51
		x"0040" & "0000011111100000", -- Address =  52
		x"0400" & "0000111111110000", -- Address =  53
		x"4000" & "0001111001111000", -- Address =  54
		x"5000" & "0011110000111100", -- Address =  55
		x"6000" & "0111100000011110", -- Address =  56
		x"1000" & "1111000000001111", -- Address =  57
		x"0100" & "1111100000011111", -- Address =  58
		x"0010" & "0111110000111110", -- Address =  59
		x"0001" & "0011111001111100", -- Address =  60
		x"0000" & "0001111111111000", -- Address =  61
		x"0000" & "0000111111110000", -- Address =  62
		x"0000" & "0000011111100000", -- Address =  63
		x"0000" & "0000111111110000", -- Address =  64
		x"0000" & "0001111111111000", -- Address =  65
		x"0000" & "0011111001111100", -- Address =  66
		x"0000" & "0111110000111110", -- Address =  67
		x"0000" & "1111100000011111", -- Address =  68
		x"0000" & "1111110000111111", -- Address =  69
		x"0000" & "0111111001111110", -- Address =  70
		x"0000" & "0011111111111100", -- Address =  71
		x"0000" & "0001111111111000", -- Address =  72
		x"0000" & "0000111111110000", -- Address =  73
		x"0000" & "0000011111100000", -- Address =  74
		x"0000" & "0000111111110000", -- Address =  75
		x"0000" & "0001111111111000", -- Address =  76
		x"0000" & "0011111111111100", -- Address =  77
		x"0000" & "0111111001111110", -- Address =  78
		x"0000" & "1111110000111111", -- Address =  79
		x"0000" & "1111111001111111", -- Address =  80
		x"0000" & "0111111111111110", -- Address =  81
		x"0000" & "0011111111111100", -- Address =  82
		x"0000" & "0001111111111000", -- Address =  83
		x"0000" & "0000111111110000", -- Address =  84
		x"0000" & "0000111111110000", -- Address =  85
		x"0000" & "0001111111111000", -- Address =  86
		x"0000" & "0011111111111100", -- Address =  87
		x"0000" & "0111111111111110", -- Address =  88
		x"0000" & "1111111111111111", -- Address =  89
		x"0000" & "0111111111111110", -- Address =  90
		x"0000" & "0011111111111100", -- Address =  91
		x"0000" & "0001111111111000", -- Address =  92
		x"0000" & "0000111111110000", -- Address =  93
		x"0000" & "0001111111111000", -- Address =  94
		x"0000" & "0011111111111100", -- Address =  95
		x"0000" & "0111111111111110", -- Address =  96
		x"0000" & "1111111111111111", -- Address =  97
		x"0000" & "0000000000000000", -- Address =  98
		x"0000" & "0000000000000000", -- Address =  99
		x"0000" & "0000000000000000", -- Address = 100
		x"0000" & "0000000000000000", -- Address = 101
		x"0000" & "0000000000000000", -- Address = 102
		x"0000" & "0000000000000000", -- Address = 103
		x"0000" & "0000000000000000", -- Address = 104
		x"0000" & "0000000000000000", -- Address = 105
		x"0000" & "0000000000000000", -- Address = 106
		x"0000" & "0000000000000000", -- Address = 107
		x"0000" & "0000000000000000", -- Address = 108
		x"0000" & "0000000000000000", -- Address = 109
		x"0000" & "0000000000000000", -- Address = 110
		x"0000" & "0000000000000000", -- Address = 111
		x"0000" & "0000000000000000", -- Address = 112
		x"0000" & "0000000000000000", -- Address = 113
		x"0000" & "0000000000000000", -- Address = 114
		x"0000" & "0000000000000000", -- Address = 115
		x"0000" & "0000000000000000", -- Address = 116
		x"0000" & "0000000000000000", -- Address = 117
		x"0000" & "0000000000000000", -- Address = 118
		x"0000" & "0000000000000000", -- Address = 119
		x"0000" & "0000000000000000", -- Address = 120
		x"0000" & "0000000000000000", -- Address = 121
		x"0000" & "0000000000000000", -- Address = 122
		x"0000" & "0000000000000000", -- Address = 123
		x"0000" & "0000000000000000", -- Address = 124
		x"0000" & "0000000000000000", -- Address = 125
		x"0000" & "0000000000000000", -- Address = 126
		x"0000" & "0000000000000000", -- Address = 127
		x"0000" & "0000000000000000", -- Address = 128
		x"0000" & "0000000000000000", -- Address = 129
		x"0000" & "0000000000000000", -- Address = 130
		x"0000" & "0000000000000000", -- Address = 131
		x"0000" & "0000000000000000", -- Address = 132
		x"0000" & "0000000000000000", -- Address = 133
		x"0000" & "0000000000000000", -- Address = 134
		x"0000" & "0000000000000000", -- Address = 135
		x"0000" & "0000000000000000", -- Address = 136
		x"0000" & "0000000000000000", -- Address = 137
		x"0000" & "0000000000000000", -- Address = 138
		x"0000" & "0000000000000000", -- Address = 139
		x"0000" & "0000000000000000", -- Address = 140
		x"0000" & "0000000000000000", -- Address = 141
		x"0000" & "0000000000000000", -- Address = 142
		x"0000" & "0000000000000000", -- Address = 143
		x"0000" & "0000000000000000", -- Address = 144
		x"0000" & "0000000000000000", -- Address = 145
		x"0000" & "0000000000000000", -- Address = 146
		x"0000" & "0000000000000000", -- Address = 147
		x"0000" & "0000000000000000", -- Address = 148
		x"0000" & "0000000000000000", -- Address = 149
		x"0000" & "0000000000000000", -- Address = 150
		x"0000" & "0000000000000000", -- Address = 151
		x"0000" & "0000000000000000", -- Address = 152
		x"0000" & "0000000000000000", -- Address = 153
		x"0000" & "0000000000000000", -- Address = 154
		x"0000" & "0000000000000000", -- Address = 155
		x"0000" & "0000000000000000", -- Address = 156
		x"0000" & "0000000000000000", -- Address = 157
		x"0000" & "0000000000000000", -- Address = 158
		x"0000" & "0000000000000000", -- Address = 159
		x"0000" & "0000000000000000", -- Address = 160
		x"0000" & "0000000000000000", -- Address = 161
		x"0000" & "0000000000000000", -- Address = 162
		x"0000" & "0000000000000000", -- Address = 163
		x"0000" & "0000000000000000", -- Address = 164
		x"0000" & "0000000000000000", -- Address = 165
		x"0000" & "0000000000000000", -- Address = 166
		x"0000" & "0000000000000000", -- Address = 167
		x"0000" & "0000000000000000", -- Address = 168
		x"0000" & "0000000000000000", -- Address = 169
		x"0000" & "0000000000000000", -- Address = 170
		x"0000" & "0000000000000000", -- Address = 171
		x"0000" & "0000000000000000", -- Address = 172
		x"0000" & "0000000000000000", -- Address = 173
		x"0000" & "0000000000000000", -- Address = 174
		x"0000" & "0000000000000000", -- Address = 175
		x"0000" & "0000000000000000", -- Address = 176
		x"0000" & "0000000000000000", -- Address = 177
		x"0000" & "0000000000000000", -- Address = 178
		x"0000" & "0000000000000000", -- Address = 179
		x"0000" & "0000000000000000", -- Address = 180
		x"0000" & "0000000000000000", -- Address = 181
		x"0000" & "0000000000000000", -- Address = 182
		x"0000" & "0000000000000000", -- Address = 183
		x"0000" & "0000000000000000", -- Address = 184
		x"0000" & "0000000000000000", -- Address = 185
		x"0000" & "0000000000000000", -- Address = 186
		x"0000" & "0000000000000000", -- Address = 187
		x"0000" & "0000000000000000", -- Address = 188
		x"0000" & "0000000000000000", -- Address = 189
		x"0000" & "0000000000000000", -- Address = 190
		x"0000" & "0000000000000000", -- Address = 191
		x"0000" & "0000000000000000", -- Address = 192
		x"0000" & "0000000000000000", -- Address = 193
		x"0000" & "0000000000000000", -- Address = 194
		x"0000" & "0000000000000000", -- Address = 195
		x"0000" & "0000000000000000", -- Address = 196
		x"0000" & "0000000000000000", -- Address = 197
		x"0000" & "0000000000000000", -- Address = 198
		x"0000" & "0000000000000000", -- Address = 199
		x"0000" & "0000000000000000", -- Address = 200
		x"0000" & "0000000000000000", -- Address = 201
		x"0000" & "0000000000000000", -- Address = 202
		x"0000" & "0000000000000000", -- Address = 203
		x"0000" & "0000000000000000", -- Address = 204
		x"0000" & "0000000000000000", -- Address = 205
		x"0000" & "0000000000000000", -- Address = 206
		x"0000" & "0000000000000000", -- Address = 207
		x"0000" & "0000000000000000", -- Address = 208
		x"0000" & "0000000000000000", -- Address = 209
		x"0000" & "0000000000000000", -- Address = 210
		x"0000" & "0000000000000000", -- Address = 211
		x"0000" & "0000000000000000", -- Address = 212
		x"0000" & "0000000000000000", -- Address = 213
		x"0000" & "0000000000000000", -- Address = 214
		x"0000" & "0000000000000000", -- Address = 215
		x"0000" & "0000000000000000", -- Address = 216
		x"0000" & "0000000000000000", -- Address = 217
		x"0000" & "0000000000000000", -- Address = 218
		x"0000" & "0000000000000000", -- Address = 219
		x"0000" & "0000000000000000", -- Address = 220
		x"0000" & "0000000000000000", -- Address = 221
		x"0000" & "0000000000000000", -- Address = 222
		x"0000" & "0000000000000000", -- Address = 223
		x"0000" & "0000000000000000", -- Address = 224
		x"0000" & "0000000000000000", -- Address = 225
		x"0000" & "0000000000000000", -- Address = 226
		x"0000" & "0000000000000000", -- Address = 227
		x"0000" & "0000000000000000", -- Address = 228
		x"0000" & "0000000000000000", -- Address = 229
		x"0000" & "0000000000000000", -- Address = 230
		x"0000" & "0000000000000000", -- Address = 231
		x"0000" & "0000000000000000", -- Address = 232
		x"0000" & "0000000000000000", -- Address = 233
		x"0000" & "0000000000000000", -- Address = 234
		x"0000" & "0000000000000000", -- Address = 235
		x"0000" & "0000000000000000", -- Address = 236
		x"0000" & "0000000000000000", -- Address = 237
		x"0000" & "0000000000000000", -- Address = 238
		x"0000" & "0000000000000000", -- Address = 239
		x"0000" & "0000000000000000", -- Address = 240
		x"0000" & "0000000000000000", -- Address = 241
		x"0000" & "0000000000000000", -- Address = 242
		x"0000" & "0000000000000000", -- Address = 243
		x"0000" & "0000000000000000", -- Address = 244
		x"0000" & "0000000000000000", -- Address = 245
		x"0000" & "0000000000000000", -- Address = 246
		x"0000" & "0000000000000000", -- Address = 247
		x"0000" & "0000000000000000", -- Address = 248
		x"0000" & "0000000000000000", -- Address = 249
		x"0000" & "0000000000000000", -- Address = 250
		x"0000" & "0000000000000000", -- Address = 251
		x"0000" & "0000000000000000", -- Address = 252
		x"0000" & "0000000000000000", -- Address = 253
		x"0000" & "0000000000000000", -- Address = 254
		x"0000" & "0000000000000000"  -- Address = 255
	);

begin

    RD <= ROM(to_integer(unsigned(A(7 downto 0))));

end architecture;
